module LUT (
    input       clk,
    input [3:0] index_0,
    input [3:0] index_1,
    input [3:0] index_2,

    output reg [11:0] addr_0,
    output reg [11:0] addr_1,
    output reg [11:0] addr_2  
);

    


    
endmodule